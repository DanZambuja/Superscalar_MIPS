library IEEE; 
use IEEE.STD_LOGIC_1164.all;  
use IEEE.STD_LOGIC_ARITH.all;

entity scoreboard_control is
    port(
        clock, reset :  in  STD_LOGIC
    );
end scoreboard_control;

architecture state_machine of scoreboard_control is


begin


end;